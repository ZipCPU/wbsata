	// Verilator lint_off UNUSED
	// These defined primitives are BIG_ENDIAN.  The first byte out is on
	// the left.  The first bit out is the LSB on the right.

				// Byte 0,	Byte 1,		Byte 2,		Byte 3
				// K.3b.5b,	D.3b.5b,	D.3b.5b,	D.3b.5b
				// Z.HGF.EDCBA
	localparam	[32:0]	P_ALIGN  = { 1'b1, 8'b101_11100, 8'b010_01010, 8'b010_01010, 8'b011_11011 },
				P_CONT   = { 1'b1, 8'b011_11100, 8'b101_01010, 8'b100_11001, 8'b100_11001 },
				P_DMAT   = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b001_10110, 8'b001_10110 },
				P_EOF    = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b110_10101, 8'b110_10101 },
				P_HOLD   = { 1'b1, 8'b011_11100, 8'b101_01010, 8'b110_10101, 8'b110_10101 },
				P_HOLDA  = { 1'b1, 8'b011_11100, 8'b101_01010, 8'b100_10101, 8'b100_10101 },
				P_PMACK  = { 1'b1, 8'b011_11100, 8'b100_10101, 8'b100_10101, 8'b100_10101 },
				P_PMNAK  = { 1'b1, 8'b011_11100, 8'b100_10101, 8'b111_10101, 8'b111_10101 },
				P_PMREQ_P= { 1'b1, 8'b011_11100, 8'b101_10101, 8'b000_10111, 8'b000_10111 },
				P_PMREQ_S= { 1'b1, 8'b011_11100, 8'b100_10101, 8'b011_10101, 8'b011_10101 },
				P_R_ERR  = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b010_10110, 8'b010_10110 },
				P_R_IP   = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b010_10101, 8'b010_10101 },
				P_R_OK   = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b001_10101, 8'b001_10101 },
				P_R_RDY  = { 1'b1, 8'b011_11100, 8'b100_10101, 8'b010_01010, 8'b010_01010 },
				P_SOF    = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b001_10111, 8'b001_10111 },
				P_SYNC   = { 1'b1, 8'b011_11100, 8'b100_10101, 8'b101_10101, 8'b101_10101 },
				P_WTRM   = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b010_11000, 8'b010_11000 },
				P_X_RDY  = { 1'b1, 8'b011_11100, 8'b101_10101, 8'b010_10111, 8'b010_10111 };
	// Verilator lint_on  UNUSED
